`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:17:05 09/01/2023 
// Design Name: 
// Module Name:    SMIX 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SMIX(
    input [31:0] word_in,
    input [1:0] index,
    input last_round,
    output [31:0] cipher_out
    );


endmodule
